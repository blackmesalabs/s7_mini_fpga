module time_stamp
(
  output wire [31:0]  time_dout
);
  assign time_dout  = 32'h5b310f03;
// Mon Jun 25 08:49:23 2018
endmodule
